`include "mux32to1_1bit.v"

module Mux32to1_32bit(input[31:0] in0, input[31:0] in1, input[31:0] in2, input[31:0] in3, input[31:0] in4, input[31:0] in5, input[31:0] in6, input[31:0] in7,
    input[31:0] in8, input[31:0] in9, input[31:0] in10, input[31:0] in11, input[31:0] in12, input[31:0] in13, input[31:0] in14, input[31:0] in15,
    input[31:0] in16, input[31:0] in17, input[31:0] in18, input[31:0] in19, input[31:0] in20, input[31:0] in21, input[31:0] in22, input[31:0] in23,
    input[31:0] in24, input[31:0] in25, input[31:0] in26, input[31:0] in27, input[31:0] in28, input[31:0] in29, input[31:0] in30, input[31:0] in31,input[4:0] select,output wire[31:0] muxOut);
   
   //WRITE YOUR CODE HERE
	Mux32to1_1bit m0(in0[0],in1[0],in2[0],in3[0],in4[0],in5[0],in6[0],in7[0],in8[0],in9[0],in10[0],in11[0],in12[0],in13[0],in14[0],in15[0],in16[0],in17[0],in18[0],in19[0],in20[0],in21[0],in22[0],in23[0],in24[0],in25[0],in26[0],in27[0],in28[0],in29[0],in30[0],in31[0], select, muxOut[0]);
    Mux32to1_1bit m1(in0[1],in1[1],in2[1],in3[1],in4[1],in5[1],in6[1],in7[1],in8[1],in9[1],in10[1],in11[1],in12[1],in13[1],in14[1],in15[1],in16[1],in17[1],in18[1],in19[1],in20[1],in21[1],in22[1],in23[1],in24[1],in25[1],in26[1],in27[1],in28[1],in29[1],in30[1],in31[1], select, muxOut[1]);
    Mux32to1_1bit m2(in0[2],in1[2],in2[2],in3[2],in4[2],in5[2],in6[2],in7[2],in8[2],in9[2],in10[2],in11[2],in12[2],in13[2],in14[2],in15[2],in16[2],in17[2],in18[2],in19[2],in20[2],in21[2],in22[2],in23[2],in24[2],in25[2],in26[2],in27[2],in28[2],in29[2],in30[2],in31[2], select, muxOut[2]);
    Mux32to1_1bit m3(in0[3],in1[3],in2[3],in3[3],in4[3],in5[3],in6[3],in7[3],in8[3],in9[3],in10[3],in11[3],in12[3],in13[3],in14[3],in15[3],in16[3],in17[3],in18[3],in19[3],in20[3],in21[3],in22[3],in23[3],in24[3],in25[3],in26[3],in27[3],in28[3],in29[3],in30[3],in31[3], select, muxOut[3]);
    Mux32to1_1bit m4(in0[4],in1[4],in2[4],in3[4],in4[4],in5[4],in6[4],in7[4],in8[4],in9[4],in10[4],in11[4],in12[4],in13[4],in14[4],in15[4],in16[4],in17[4],in18[4],in19[4],in20[4],in21[4],in22[4],in23[4],in24[4],in25[4],in26[4],in27[4],in28[4],in29[4],in30[4],in31[4], select, muxOut[4]);
    Mux32to1_1bit m5(in0[5],in1[5],in2[5],in3[5],in4[5],in5[5],in6[5],in7[5],in8[5],in9[5],in10[5],in11[5],in12[5],in13[5],in14[5],in15[5],in16[5],in17[5],in18[5],in19[5],in20[5],in21[5],in22[5],in23[5],in24[5],in25[5],in26[5],in27[5],in28[5],in29[5],in30[5],in31[5], select, muxOut[5]);
    Mux32to1_1bit m6(in0[6],in1[6],in2[6],in3[6],in4[6],in5[6],in6[6],in7[6],in8[6],in9[6],in10[6],in11[6],in12[6],in13[6],in14[6],in15[6],in16[6],in17[6],in18[6],in19[6],in20[6],in21[6],in22[6],in23[6],in24[6],in25[6],in26[6],in27[6],in28[6],in29[6],in30[6],in31[6], select, muxOut[6]);
    Mux32to1_1bit m7(in0[7],in1[7],in2[7],in3[7],in4[7],in5[7],in6[7],in7[7],in8[7],in9[7],in10[7],in11[7],in12[7],in13[7],in14[7],in15[7],in16[7],in17[7],in18[7],in19[7],in20[7],in21[7],in22[7],in23[7],in24[7],in25[7],in26[7],in27[7],in28[7],in29[7],in30[7],in31[7], select, muxOut[7]);
    Mux32to1_1bit m8(in0[8],in1[8],in2[8],in3[8],in4[8],in5[8],in6[8],in7[8],in8[8],in9[8],in10[8],in11[8],in12[8],in13[8],in14[8],in15[8],in16[8],in17[8],in18[8],in19[8],in20[8],in21[8],in22[8],in23[8],in24[8],in25[8],in26[8],in27[8],in28[8],in29[8],in30[8],in31[8], select, muxOut[8]);
    Mux32to1_1bit m9(in0[9],in1[9],in2[9],in3[9],in4[9],in5[9],in6[9],in7[9],in8[9],in9[9],in10[9],in11[9],in12[9],in13[9],in14[9],in15[9],in16[9],in17[9],in18[9],in19[9],in20[9],in21[9],in22[9],in23[9],in24[9],in25[9],in26[9],in27[9],in28[9],in29[9],in30[9],in31[9], select, muxOut[9]);
    Mux32to1_1bit m10(in0[10],in1[10],in2[10],in3[10],in4[10],in5[10],in6[10],in7[10],in8[10],in9[10],in10[10],in11[10],in12[10],in13[10],in14[10],in15[10],in16[10],in17[10],in18[10],in19[10],in20[10],in21[10],in22[10],in23[10],in24[10],in25[10],in26[10],in27[10],in28[10],in29[10],in30[10],in31[10], select, muxOut[10]);
    Mux32to1_1bit m11(in0[11],in1[11],in2[11],in3[11],in4[11],in5[11],in6[11],in7[11],in8[11],in9[11],in10[11],in11[11],in12[11],in13[11],in14[11],in15[11],in16[11],in17[11],in18[11],in19[11],in20[11],in21[11],in22[11],in23[11],in24[11],in25[11],in26[11],in27[11],in28[11],in29[11],in30[11],in31[11], select, muxOut[11]);
    Mux32to1_1bit m12(in0[12],in1[12],in2[12],in3[12],in4[12],in5[12],in6[12],in7[12],in8[12],in9[12],in10[12],in11[12],in12[12],in13[12],in14[12],in15[12],in16[12],in17[12],in18[12],in19[12],in20[12],in21[12],in22[12],in23[12],in24[12],in25[12],in26[12],in27[12],in28[12],in29[12],in30[12],in31[12], select, muxOut[12]);
    Mux32to1_1bit m13(in0[13],in1[13],in2[13],in3[13],in4[13],in5[13],in6[13],in7[13],in8[13],in9[13],in10[13],in11[13],in12[13],in13[13],in14[13],in15[13],in16[13],in17[13],in18[13],in19[13],in20[13],in21[13],in22[13],in23[13],in24[13],in25[13],in26[13],in27[13],in28[13],in29[13],in30[13],in31[13], select, muxOut[13]);
    Mux32to1_1bit m14(in0[14],in1[14],in2[14],in3[14],in4[14],in5[14],in6[14],in7[14],in8[14],in9[14],in10[14],in11[14],in12[14],in13[14],in14[14],in15[14],in16[14],in17[14],in18[14],in19[14],in20[14],in21[14],in22[14],in23[14],in24[14],in25[14],in26[14],in27[14],in28[14],in29[14],in30[14],in31[14], select, muxOut[14]);
    Mux32to1_1bit m15(in0[15],in1[15],in2[15],in3[15],in4[15],in5[15],in6[15],in7[15],in8[15],in9[15],in10[15],in11[15],in12[15],in13[15],in14[15],in15[15],in16[15],in17[15],in18[15],in19[15],in20[15],in21[15],in22[15],in23[15],in24[15],in25[15],in26[15],in27[15],in28[15],in29[15],in30[15],in31[15], select, muxOut[15]);
    Mux32to1_1bit m16(in0[16],in1[16],in2[16],in3[16],in4[16],in5[16],in6[16],in7[16],in8[16],in9[16],in10[16],in11[16],in12[16],in13[16],in14[16],in15[16],in16[16],in17[16],in18[16],in19[16],in20[16],in21[16],in22[16],in23[16],in24[16],in25[16],in26[16],in27[16],in28[16],in29[16],in30[16],in31[16], select, muxOut[16]);
    Mux32to1_1bit m17(in0[17],in1[17],in2[17],in3[17],in4[17],in5[17],in6[17],in7[17],in8[17],in9[17],in10[17],in11[17],in12[17],in13[17],in14[17],in15[17],in16[17],in17[17],in18[17],in19[17],in20[17],in21[17],in22[17],in23[17],in24[17],in25[17],in26[17],in27[17],in28[17],in29[17],in30[17],in31[17], select, muxOut[17]);
    Mux32to1_1bit m18(in0[18],in1[18],in2[18],in3[18],in4[18],in5[18],in6[18],in7[18],in8[18],in9[18],in10[18],in11[18],in12[18],in13[18],in14[18],in15[18],in16[18],in17[18],in18[18],in19[18],in20[18],in21[18],in22[18],in23[18],in24[18],in25[18],in26[18],in27[18],in28[18],in29[18],in30[18],in31[18], select, muxOut[18]);
    Mux32to1_1bit m19(in0[19],in1[19],in2[19],in3[19],in4[19],in5[19],in6[19],in7[19],in8[19],in9[19],in10[19],in11[19],in12[19],in13[19],in14[19],in15[19],in16[19],in17[19],in18[19],in19[19],in20[19],in21[19],in22[19],in23[19],in24[19],in25[19],in26[19],in27[19],in28[19],in29[19],in30[19],in31[19], select, muxOut[19]);
    Mux32to1_1bit m20(in0[20],in1[20],in2[20],in3[20],in4[20],in5[20],in6[20],in7[20],in8[20],in9[20],in10[20],in11[20],in12[20],in13[20],in14[20],in15[20],in16[20],in17[20],in18[20],in19[20],in20[20],in21[20],in22[20],in23[20],in24[20],in25[20],in26[20],in27[20],in28[20],in29[20],in30[20],in31[20], select, muxOut[20]);
    Mux32to1_1bit m21(in0[21],in1[21],in2[21],in3[21],in4[21],in5[21],in6[21],in7[21],in8[21],in9[21],in10[21],in11[21],in12[21],in13[21],in14[21],in15[21],in16[21],in17[21],in18[21],in19[21],in20[21],in21[21],in22[21],in23[21],in24[21],in25[21],in26[21],in27[21],in28[21],in29[21],in30[21],in31[21], select, muxOut[21]);
    Mux32to1_1bit m22(in0[22],in1[22],in2[22],in3[22],in4[22],in5[22],in6[22],in7[22],in8[22],in9[22],in10[22],in11[22],in12[22],in13[22],in14[22],in15[22],in16[22],in17[22],in18[22],in19[22],in20[22],in21[22],in22[22],in23[22],in24[22],in25[22],in26[22],in27[22],in28[22],in29[22],in30[22],in31[22], select, muxOut[22]);
    Mux32to1_1bit m23(in0[23],in1[23],in2[23],in3[23],in4[23],in5[23],in6[23],in7[23],in8[23],in9[23],in10[23],in11[23],in12[23],in13[23],in14[23],in15[23],in16[23],in17[23],in18[23],in19[23],in20[23],in21[23],in22[23],in23[23],in24[23],in25[23],in26[23],in27[23],in28[23],in29[23],in30[23],in31[23], select, muxOut[23]);
    Mux32to1_1bit m24(in0[24],in1[24],in2[24],in3[24],in4[24],in5[24],in6[24],in7[24],in8[24],in9[24],in10[24],in11[24],in12[24],in13[24],in14[24],in15[24],in16[24],in17[24],in18[24],in19[24],in20[24],in21[24],in22[24],in23[24],in24[24],in25[24],in26[24],in27[24],in28[24],in29[24],in30[24],in31[24], select, muxOut[24]);
    Mux32to1_1bit m25(in0[25],in1[25],in2[25],in3[25],in4[25],in5[25],in6[25],in7[25],in8[25],in9[25],in10[25],in11[25],in12[25],in13[25],in14[25],in15[25],in16[25],in17[25],in18[25],in19[25],in20[25],in21[25],in22[25],in23[25],in24[25],in25[25],in26[25],in27[25],in28[25],in29[25],in30[25],in31[25], select, muxOut[25]);
    Mux32to1_1bit m26(in0[26],in1[26],in2[26],in3[26],in4[26],in5[26],in6[26],in7[26],in8[26],in9[26],in10[26],in11[26],in12[26],in13[26],in14[26],in15[26],in16[26],in17[26],in18[26],in19[26],in20[26],in21[26],in22[26],in23[26],in24[26],in25[26],in26[26],in27[26],in28[26],in29[26],in30[26],in31[26], select, muxOut[26]);
    Mux32to1_1bit m27(in0[27],in1[27],in2[27],in3[27],in4[27],in5[27],in6[27],in7[27],in8[27],in9[27],in10[27],in11[27],in12[27],in13[27],in14[27],in15[27],in16[27],in17[27],in18[27],in19[27],in20[27],in21[27],in22[27],in23[27],in24[27],in25[27],in26[27],in27[27],in28[27],in29[27],in30[27],in31[27], select, muxOut[27]);
    Mux32to1_1bit m28(in0[28],in1[28],in2[28],in3[28],in4[28],in5[28],in6[28],in7[28],in8[28],in9[28],in10[28],in11[28],in12[28],in13[28],in14[28],in15[28],in16[28],in17[28],in18[28],in19[28],in20[28],in21[28],in22[28],in23[28],in24[28],in25[28],in26[28],in27[28],in28[28],in29[28],in30[28],in31[28], select, muxOut[28]);
    Mux32to1_1bit m29(in0[29],in1[29],in2[29],in3[29],in4[29],in5[29],in6[29],in7[29],in8[29],in9[29],in10[29],in11[29],in12[29],in13[29],in14[29],in15[29],in16[29],in17[29],in18[29],in19[29],in20[29],in21[29],in22[29],in23[29],in24[29],in25[29],in26[29],in27[29],in28[29],in29[29],in30[29],in31[29], select, muxOut[29]);
    Mux32to1_1bit m30(in0[30],in1[30],in2[30],in3[30],in4[30],in5[30],in6[30],in7[30],in8[30],in9[30],in10[30],in11[30],in12[30],in13[30],in14[30],in15[30],in16[30],in17[30],in18[30],in19[30],in20[30],in21[30],in22[30],in23[30],in24[30],in25[30],in26[30],in27[30],in28[30],in29[30],in30[30],in31[30], select, muxOut[30]);
    Mux32to1_1bit m31(in0[31],in1[31],in2[31],in3[31],in4[31],in5[31],in6[31],in7[31],in8[31],in9[31],in10[31],in11[31],in12[31],in13[31],in14[31],in15[31],in16[31],in17[31],in18[31],in19[31],in20[31],in21[31],in22[31],in23[31],in24[31],in25[31],in26[31],in27[31],in28[31],in29[31],in30[31],in31[31], select, muxOut[31]);


endmodule
